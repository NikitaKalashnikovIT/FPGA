test 1 br1
